library verilog;
use verilog.vl_types.all;
entity relogio_vlg_sample_tst is
    port(
        clockIn         : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end relogio_vlg_sample_tst;

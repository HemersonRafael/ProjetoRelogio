--library ieee;
--
--use ieee.std_logic_1164.all;
--
--entity convesorBD is
--	port(vectorBits: std_logic (5 downto 0));
--	
--end convesorBD;
--
--architecture hardware of convesorBD is
--signal soma : integer := 0;
--soma <= to_integer(unsigned(vectorBits));
--end hardware;
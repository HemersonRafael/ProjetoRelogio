library verilog;
use verilog.vl_types.all;
entity contadorHMS_vlg_vec_tst is
end contadorHMS_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity contadorCrescente_vlg_vec_tst is
end contadorCrescente_vlg_vec_tst;
